package RISCV_CORE_CONFIG_BENCH is
	constant PERIOD : time := 20 ns;
	constant HALF_PERIOD : time := PERIOD / 2;
	constant QUARTER_PERIOD : time := PERIOD / 4;
end package RISCV_CORE_CONFIG_BENCH;
